module secondInterval_zgrankin(clock, reset, );
	input clock;
	input reset;
	
	assign out = (count == 25'd24999999)

	if (count == 25'd24999999)
		count = 25'd0;